
module sys (
	clk_clk,
	master_0_master_reset_reset,
	pio_0_external_connection_export,
	reset_reset_n);	

	input		clk_clk;
	output		master_0_master_reset_reset;
	output	[7:0]	pio_0_external_connection_export;
	input		reset_reset_n;
endmodule
