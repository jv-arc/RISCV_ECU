// Debug values for the convention used in the C code for flags

parameter NORMAL = 8'h00;
parameter SUCCESS = 8'hF0;
parameter FAILURE = 8'hFF;

parameter MAIN = 8'h00;
parameter WHILE = 8'h01;
parameter FUNC = 8'h02;
parameter SETUP = 8'h03;
parameter ISR = 8'h04;
