
module sys (
	clk_clk,
	gpio_a_dir_external_connection_export,
	gpio_a_r_external_connection_export,
	gpio_a_w_external_connection_export,
	gpio_b_dir_external_connection_export,
	gpio_b_r_external_connection_export,
	gpio_b_w_external_connection_export,
	master_0_master_reset_reset,
	pio_r_one_external_connection_export,
	pio_w_one_external_connection_export,
	pio_w_two_external_connection_export,
	pulpino_0_config_testmode_i,
	pulpino_0_config_fetch_enable_i,
	pulpino_0_config_clock_gating_i,
	pulpino_0_config_boot_addr_i,
	reset_reset_n);	

	input		clk_clk;
	output	[31:0]	gpio_a_dir_external_connection_export;
	input	[31:0]	gpio_a_r_external_connection_export;
	output	[31:0]	gpio_a_w_external_connection_export;
	output	[31:0]	gpio_b_dir_external_connection_export;
	input	[31:0]	gpio_b_r_external_connection_export;
	output	[31:0]	gpio_b_w_external_connection_export;
	output		master_0_master_reset_reset;
	input	[31:0]	pio_r_one_external_connection_export;
	output	[31:0]	pio_w_one_external_connection_export;
	output	[31:0]	pio_w_two_external_connection_export;
	input		pulpino_0_config_testmode_i;
	input		pulpino_0_config_fetch_enable_i;
	input		pulpino_0_config_clock_gating_i;
	input	[31:0]	pulpino_0_config_boot_addr_i;
	input		reset_reset_n;
endmodule
